/* ==================================================
 * Filename: %FFILE% 
 * Date    : %DATE%
 * Author  : %USER%
 * Contact : %MAIL%
 * ==================================================
 */

%HERE%
